/*
1. The role of the "sequencer" is to initiate the "sequence"
2. Sequencer can send item ("item" is created by sequence) to the driver
*/

typedef uvm_sequencer #(my_transaction) my_sequencer;
