typedef uvm_sequencer #(my_seq_item) CompSeqr;
