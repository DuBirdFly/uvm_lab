module router_iport (
    input                   clk,
    input                   reset_n,

    input                   i_frame,
    input                   i_data,
    output                  o_dst_addr,

    input                   i_gnt,
    output                  o_req

);
















endmodule