typedef uvm_sequencer #(TrAxi) AxiMasterSeqr;