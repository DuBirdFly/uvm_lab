typedef uvm_sequencer #(TrApb) ApbMasterSeqr;