module router_iport (
    input                   clk,
    input                   reset_n,

    input                   i_frame,
    input                   i_valid,
    input                   i_data,

    output                  o_req,
    output                  o_data

);



endmodule