class CfgAgt extend uvm_object;

    /* 声明变量 */
    uvm_active_passive_enum is_active = UVM_ACTIVE;
    int unsigned pad_cycle = 5;
    virtual IntfDut intf_dut;

    /* 注册变量 */












endclass