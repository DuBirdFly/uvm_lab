typedef uvm_sequencer #(TrApb) SeqrApb;