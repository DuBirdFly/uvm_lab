typedef uvm_sequencer #(MySeqItem) CompSeqr;
