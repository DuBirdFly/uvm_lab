`define APB_WIDTH 32
`define APB_DEPTH 16
